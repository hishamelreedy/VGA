//Verilog HDL for "cuaic", "not" "functional"


module not1  ( input wire x, output wire y);
assign y=~x;
endmodule
